default.vhd#16096#0#0#{0000}>-{0000}